// femtorv32, a minimalistic RISC-V RV32I core
//    (minus SYSTEM and FENCE that are not implemented)
//
//       Bruno Levy, 2020-2021
//
// This file: FGA: Femto Graphics Adapter
//   Note: VRAM is write-only ! (the read port is used by HDMI)
//   Mode 1: 320x200x16bpp. 

`include "HDMI_clock.v"
`include "TMDS_encoder.v"

module FGA(
    input wire 	      clk,         // system clock
    input wire 	      sel,         // if zero, writes are ignored
    input wire [3:0]  mem_wmask,   // mem write mask and strobe /write Legal values are 000,0001,0010,0100,1000,0011,1100,1111	   
    input wire [16:0] mem_address, // address in graphic memory (128K), word-aligned
    input wire [31:0] mem_wdata,   // data to be written

    input wire        pixel_clk,   // 25 MHz	   
    output wire [3:0] gpdi_dp      // HDMI signals, blue, green, red, clock
                                   // dgpi_dn generated by pins (see ulx3s.lpf)
);

   wire [14:0] vram_word_address = mem_address[16:2];

   reg [31:0] VRAM[32767:0];

   // write VRAM (interface with processor)
   always @(posedge clk) begin
      if(sel) begin
	 if(mem_wmask[0]) VRAM[vram_word_address][ 7:0 ] <= mem_wdata[ 7:0 ];
	 if(mem_wmask[1]) VRAM[vram_word_address][15:8 ] <= mem_wdata[15:8 ];
	 if(mem_wmask[2]) VRAM[vram_word_address][23:16] <= mem_wdata[23:16];
	 if(mem_wmask[3]) VRAM[vram_word_address][31:24] <= mem_wdata[31:24];	 
      end 
   end

   /************************* HDMI signal generation ***************************/
   
   // This part is just like a VGA generator.
   reg [9:0] X, Y;   // current pixel coordinates
   reg hSync, vSync; // horizontal and vertical synchronization
   reg DrawArea;     // asserted if current pixel is in drawing area
   always @(posedge pixel_clk) begin
      DrawArea <= (X<640) && (Y<480);
      X <= (X==799) ? 0 : X+1;
      if(X==799) Y <= (Y==524) ? 0 : Y+1;
      hSync <= (X>=656) && (X<752);
      vSync <= (Y>=490) && (Y<492);
   end

   // Fetch pixel data
   reg [16:0] pix_address;
   reg [16:0] row_start;
   reg [15:0] pix_data;
   always @(posedge pixel_clk) begin
      if(X == 0) begin
	 if(Y == 0) begin
	    row_start   <= 0;
	    pix_address <= 0;
	 end else begin
	    if(Y[0]) begin
	       row_start <= row_start + 640;
	       pix_address <= row_start + 640;
	    end else begin
	       pix_address <= row_start;	       
	    end
	 end
      end 
      // Increment pix_address every 4 X (2 because 320x200->640x400 and 2 because 16 bpp)
      if(X[1:0] == 2'b11) pix_address <= pix_address + 4;

      // Draw 640x400 zone, and hide first pixel row (fetch delay)      
      // Select word's 16msb or 16lsbs based on X[1] (again, every 4 X)
      pix_data <=  (X == 0 || Y > 400) ? 0 : 
		   X[1] ? VRAM[pix_address[16:2]][31:16] : VRAM[pix_address[16:2]][15:0];
   end
   
   // Decode pixel data:  RRRRR GGGGG 0 BBBBB
   wire [7:0] R = {pix_data[15:11],3'b000};
   wire [7:0] G = {pix_data[10:5], 2'b00 };
   wire [7:0] B = {pix_data[4:0],  3'b000};

   // RGB TMDS encoding
   // Generate 10-bits TMDS red,green,blue signals. Blue embeds HSync/VSync in its 
   // control part.
   //
   // Note: Yosys finds a combinatorial loop here, but I do not understand why (and
   // it seems to work though). TO BE UNDERSTOOD.
   wire [9:0] TMDS_R, TMDS_G, TMDS_B;
   TMDS_encoder encode_R(.clk(pixel_clk), .VD(R), .CD(2'b00)        , .VDE(DrawArea), .TMDS(TMDS_R));
   TMDS_encoder encode_G(.clk(pixel_clk), .VD(G), .CD(2'b00)        , .VDE(DrawArea), .TMDS(TMDS_G));
   TMDS_encoder encode_B(.clk(pixel_clk), .VD(B), .CD({vSync,hSync}), .VDE(DrawArea), .TMDS(TMDS_B));

   // 250 MHz clock 
   // This one needs some FPGA-specific specialized blocks (a PLL).
   wire clk_TMDS; // The 250 MHz clock used by the serializers.
   HDMI_clock hdmi_clock(.clk(pixel_clk), .hdmi_clk(clk_TMDS));

   // Modulo-10 clock divider
   reg [9:0] TMDS_mod10=1;
   wire      TMDS_shift_load = TMDS_mod10[9];
   always @(posedge clk_TMDS) TMDS_mod10 <= {TMDS_mod10[8:0],TMDS_mod10[9]};

   // Shifters
   // Every 10 clocks, we get a fresh R,G,B triplet from the TMDS encoders,
   // else we shift.
   reg [9:0] TMDS_shift_R=0, TMDS_shift_G=0, TMDS_shift_B=0;
   always @(posedge clk_TMDS) begin
      TMDS_shift_R <= TMDS_shift_load ? TMDS_R : {1'b0,TMDS_shift_R[9:1]};
      TMDS_shift_G <= TMDS_shift_load ? TMDS_G : {1'b0,TMDS_shift_G[9:1]};
      TMDS_shift_B <= TMDS_shift_load ? TMDS_B : {1'b0,TMDS_shift_B[9:1]};	
   end

   // HDMI signal, positive part of the differential pairs
   // (negative part generated by the pins, see ulx3s.lpf)
   assign gpdi_dp[2] = TMDS_shift_R[0];
   assign gpdi_dp[1] = TMDS_shift_G[0];
   assign gpdi_dp[0] = TMDS_shift_B[0];
   assign gpdi_dp[3] = pixel_clk;

endmodule
	   
