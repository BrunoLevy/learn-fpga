// femtorv32, a minimalistic RISC-V RV32I core
//       Bruno Levy, 2020-2021
//
// This file: FGA: Femto Graphics Adapter
//   Note: VRAM is write-only ! (the read port is used by HDMI)
//   Mode 1: 320x200x16bpp. 

`include "HDMI_clock.v"
`include "TMDS_encoder.v"

module FGA(
    input wire 	      clk,         // system clock
    input wire 	      sel,         // if zero, writes are ignored
    input wire [3:0]  mem_wmask,   // mem write mask and strobe
    input wire [16:0] mem_address, // address in graphic memory (128K), word-aligned
    input wire [31:0] mem_wdata,   // data to be written

    input wire        pixel_clk,   // 25 MHz	   
    output wire [3:0] gpdi_dp,     // HDMI signals, blue, green, red, clock
                                   // dgpi_dn generated by pins (see ulx3s.lpf)

    input  wire io_wstrb,
    input  wire io_rstrb,
    input  wire sel_cntl,          // select control register (R/W)
    input  wire sel_dat,           // select data in (W)
    output wire	[31:0] rdata       // data read from register
);

   reg [31:0] VRAM[32767:0];
   reg [23:0] PALETTE[255:0];
   reg [1:0]  MODE;
   reg [14:0] ORIGIN;

   /************************* HDMI signal generation ***************************/

   localparam MODE_320x200x16bpp = 2'b00;
   localparam MODE_320x200x8bpp  = 2'b01;
   localparam MODE_640x400x4bpp  = 2'b10;
   
   // This part is just like a VGA generator.
   reg  [9:0] X, Y;   // current pixel coordinates
   reg hSync, vSync; // horizontal and vertical synchronization
   reg DrawArea;     // asserted if current pixel is in drawing area
   reg mem_busy;     // asserted if memory transfer is running.
   
   // read control register
   assign rdata = (io_rstrb && sel_cntl) ? 
                  {(Y >= 400),(X >= 640),DrawArea,mem_busy,4'b0,2'b0,X,2'b0,Y} : 
                  32'b0;
   
   always @(posedge pixel_clk) begin
      DrawArea <= (X<640) && (Y<480);
      X        <= (X==799) ? 0 : X+1;
      if(X==799) Y <= (Y==524) ? 0 : Y+1;
      hSync <= (X>=656) && (X<752);
      vSync <= (Y>=490) && (Y<492);
   end

   reg [14:0] pix_word_address;
   reg [14:0] row_start_word_address;
   reg [15:0] pix_data;
   reg [7:0]  R,G,B;

   always @(posedge pixel_clk) begin
      case(MODE)
	
	MODE_320x200x16bpp: begin
	   if(X == 0) begin
	      if(Y == 0) begin
		 row_start_word_address <= ORIGIN;
		 pix_word_address       <= ORIGIN;
	      end else begin
		 // Increment row address every 2 Y (2 because 320x200->640x400)
		 if(Y[0]) begin
		    row_start_word_address <= row_start_word_address + 320*2/4;
		    pix_word_address       <= row_start_word_address + 320*2/4;
		 end else begin
		    pix_word_address <= row_start_word_address;	       
		 end
	      end
	   end 
	   
	   if(X[1:0] == 2'b11) pix_word_address <= pix_word_address + 1;
	   
	   // Select word's 16msb or 16lsbs based on X[1] (again, every 4 X)
	   if(X[1]) begin 
	      R <= {VRAM[pix_word_address][31:27],3'b000};
	      G <= {VRAM[pix_word_address][26:21],2'b00 };
	      B <= {VRAM[pix_word_address][20:16],3'b000};
	   end else begin
	      R <= {VRAM[pix_word_address][15:11],3'b000};
	      G <= {VRAM[pix_word_address][10:5 ],2'b00 };
	      B <= {VRAM[pix_word_address][ 4:0 ],3'b000};
	   end
	   
	   // First pixel is boring, normally I should prefetch it...
	   if(X == 0 || Y >= 400) begin R <= 0; G <= 0; B <= 0; end
	end
	MODE_320x200x8bpp: begin
	end
	MODE_640x400x4bpp: begin
	end
      endcase
   end
   
   // RGB TMDS encoding
   // Generate 10-bits TMDS red,green,blue signals. Blue embeds HSync/VSync in its 
   // control part.
   wire [9:0] TMDS_R, TMDS_G, TMDS_B;
   TMDS_encoder encode_R(.clk(pixel_clk), .VD(R), .CD(2'b00)        , .VDE(DrawArea), .TMDS(TMDS_R));
   TMDS_encoder encode_G(.clk(pixel_clk), .VD(G), .CD(2'b00)        , .VDE(DrawArea), .TMDS(TMDS_G));
   TMDS_encoder encode_B(.clk(pixel_clk), .VD(B), .CD({vSync,hSync}), .VDE(DrawArea), .TMDS(TMDS_B));

   // 250 MHz clock 
   // This one needs some FPGA-specific specialized blocks (a PLL).
   wire clk_TMDS; // The 250 MHz clock used by the serializers.
   HDMI_clock hdmi_clock(.clk(pixel_clk), .hdmi_clk(clk_TMDS));

   // Modulo-10 clock divider (my version, using a 1-hot in a 10 bits ring)
   reg [9:0] TMDS_mod10=1;
   wire      TMDS_shift_load = TMDS_mod10[9];
   always @(posedge clk_TMDS) TMDS_mod10 <= {TMDS_mod10[8:0],TMDS_mod10[9]};

   // Shifters
   // Every 10 clocks, we get a fresh R,G,B triplet from the TMDS encoders,
   // else we shift.
   reg [9:0] TMDS_shift_R=0, TMDS_shift_G=0, TMDS_shift_B=0;
   always @(posedge clk_TMDS) begin
      TMDS_shift_R <= TMDS_shift_load ? TMDS_R : {1'b0,TMDS_shift_R[9:1]};
      TMDS_shift_G <= TMDS_shift_load ? TMDS_G : {1'b0,TMDS_shift_G[9:1]};
      TMDS_shift_B <= TMDS_shift_load ? TMDS_B : {1'b0,TMDS_shift_B[9:1]};	
   end

   // HDMI signal, positive part of the differential pairs
   // (negative part generated by the pins, see ulx3s.lpf)
   assign gpdi_dp[2] = TMDS_shift_R[0];
   assign gpdi_dp[1] = TMDS_shift_G[0];
   assign gpdi_dp[0] = TMDS_shift_B[0];
   assign gpdi_dp[3] = pixel_clk;

   /*************************************************************************/

   // control register - commands

   localparam SET_MODE       = 8'd0; 
   localparam SET_PALETTE_R  = 8'd1; 
   localparam SET_PALETTE_G  = 8'd2; 
   localparam SET_PALETTE_B  = 8'd3; 
   localparam SET_WWINDOW_X  = 8'd4;
   localparam SET_WWINDOW_Y  = 8'd5;
   localparam SET_ORIGIN     = 8'd6;
   
   
   // Emulation of SSD1351 OLED display.
   // - write window command, two commands:
   //     (send 32 bits to IO_FGA_CNTL hardware register)
   //   CMD=4: SET_WWINDOW_X: X2[11:0] X1[11:0] CMD[7:0]
   //   CMD=5: SET_WWINDOW_Y: Y2[11:0] Y1[11:0] CMD[7:0]
   //
   // - write data: send 8 bits to IO_FGA_DAT hardware register
   //    MSB first, encoding follows SSD1351: RRRRR GGGGG 0 BBBBB
   
   reg[11:0] window_x1, window_x2, window_y1, window_y2, window_x, window_y;
   reg[15:0] window_row_start;
   reg[15:0] window_hword_address;   
   
   always @(posedge clk) begin
      if(io_wstrb) begin
	 if(sel_cntl) begin
	    /* verilator lint_off CASEINCOMPLETE */
	    case(mem_wdata[7:0])
	      SET_MODE:      MODE <= mem_wdata[1:0];
	      SET_ORIGIN:    ORIGIN <= mem_wdata[16:2]; // the two LSBs are ignored
	      SET_PALETTE_R: PALETTE[mem_wdata[15:8]][7:0]   <= mem_wdata[23:16];
	      SET_PALETTE_G: PALETTE[mem_wdata[15:8]][15:8]  <= mem_wdata[23:16];
	      SET_PALETTE_B: PALETTE[mem_wdata[15:8]][23:16] <= mem_wdata[23:16];
	      SET_WWINDOW_X: begin 
		 window_x1 <= mem_wdata[19:8];
		 window_x2 <= mem_wdata[31:20];
		 window_x  <= mem_wdata[19:8];
		 mem_busy  <= 1'b1;
	      end
	      SET_WWINDOW_Y: begin 
		 window_y1 <= mem_wdata[19:8];
		 window_y2 <= mem_wdata[31:20];
		 window_y  <= mem_wdata[19:8];
		 mem_busy  <= 1'b1;
		 /* verilator lint_off WIDTH */
		 window_row_start     <= mem_wdata[19:8] * 320 + window_x1;
		 window_hword_address <= mem_wdata[19:8] * 320 + window_x1;
		 /* verilator lint_on WIDTH */		 
	      end
	    endcase
	    /* verilator lint_on CASEINCOMPLETE */	    
	 end else if(sel_dat) begin // one byte of data sent to IO_FGA_DAT
	                            // increment pixel address.
	    window_hword_address <= window_hword_address + 1;
	    window_x             <= window_x + 1;	    
	    if(window_x == window_x2) begin
	       if(window_y == window_y2) begin
		  mem_busy <= 1'b0;
	       end else begin
	          window_y <= window_y+1;
		  window_x <= window_x1;
		  window_hword_address <= window_row_start + 320;
		  window_row_start     <= window_row_start + 320;
	       end
	    end 
         end // if (sel_dat)
      end // if (wstrb)
   end // always @ (posedge clk)

   
   // write VRAM (interface with processor)
   wire [14:0] vram_word_address = mem_address[16:2];
   always @(posedge clk) begin
      if(io_wstrb) begin
         if(sel_dat && mem_busy) begin // one byte of data sent to IO_FGA_DAT
	                               // write data to VRAM.
	    case(window_hword_address[0])
	       1'b0: VRAM[window_hword_address[15:1]][15:0 ] <= mem_wdata[15:0];
	       1'b1: VRAM[window_hword_address[15:1]][31:16] <= mem_wdata[15:0];
	    endcase
	 end
      end else if(sel && !mem_busy) begin
	 if(mem_wmask[0]) VRAM[vram_word_address][ 7:0 ] <= mem_wdata[ 7:0 ];
	 if(mem_wmask[1]) VRAM[vram_word_address][15:8 ] <= mem_wdata[15:8 ];
	 if(mem_wmask[2]) VRAM[vram_word_address][23:16] <= mem_wdata[23:16];
	 if(mem_wmask[3]) VRAM[vram_word_address][31:24] <= mem_wdata[31:24];	 
      end 
   end
   
endmodule
	   
